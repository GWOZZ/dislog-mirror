library verilog;
use verilog.vl_types.all;
entity TAREA1_A_vlg_vec_tst is
end TAREA1_A_vlg_vec_tst;
