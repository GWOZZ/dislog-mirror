library verilog;
use verilog.vl_types.all;
entity TAREA1_D is
    port(
        A1              : out    vl_logic;
        SW              : in     vl_logic_vector(2 downto 0);
        B1              : out    vl_logic;
        C1              : out    vl_logic;
        D1              : out    vl_logic;
        E1              : out    vl_logic;
        F1              : out    vl_logic;
        G1              : out    vl_logic;
        A2              : out    vl_logic;
        B2              : out    vl_logic;
        C2              : out    vl_logic;
        D2              : out    vl_logic;
        E2              : out    vl_logic;
        F2              : out    vl_logic;
        G2              : out    vl_logic
    );
end TAREA1_D;
