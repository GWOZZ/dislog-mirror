library verilog;
use verilog.vl_types.all;
entity TAREA1_A_vlg_check_tst is
    port(
        Disp            : in     vl_logic_vector(6 downto 0);
        sampler_rx      : in     vl_logic
    );
end TAREA1_A_vlg_check_tst;
