library verilog;
use verilog.vl_types.all;
entity TAREA1_A_vlg_check_tst is
    port(
        LED             : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end TAREA1_A_vlg_check_tst;
