library verilog;
use verilog.vl_types.all;
entity TAREA1_D_vlg_check_tst is
    port(
        A1              : in     vl_logic;
        A2              : in     vl_logic;
        B1              : in     vl_logic;
        B2              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        D1              : in     vl_logic;
        D2              : in     vl_logic;
        E1              : in     vl_logic;
        E2              : in     vl_logic;
        F1              : in     vl_logic;
        F2              : in     vl_logic;
        G1              : in     vl_logic;
        G2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TAREA1_D_vlg_check_tst;
