library verilog;
use verilog.vl_types.all;
entity tarea1_vlg_vec_tst is
end tarea1_vlg_vec_tst;
